netcdf simple.nc {
  dimensions:
    lon = 360;
    lat = 180;
    time = UNLIMITED;   // (31 currently)
  variables:
    double lon(lon=360);
      :standard_name = "longitude";
      :long_name = "longitude";
      :units = "degrees_east";
      :axis = "X";

    double lat(lat=180);
      :standard_name = "latitude";
      :long_name = "latitude";
      :units = "degrees_north";
      :axis = "Y";

    double time(time=31);
      :standard_name = "time";
      :units = "days since 2016-01-01 00:00:00";
      :calendar = "proleptic_gregorian";

    float p(time=31, lat=180, lon=360);
      :long_name = "first guess daily product version 1 precipitation per grid";
      :units = "mm/day";
      :code = 20; // int
      :_FillValue = -99999.99f; // float

    float sd(time=31, lat=180, lon=360);
      :long_name = "first guess daily product version 1 standard deviation per grid";
      :units = "mm/day";
      :code = 22; // int
      :_FillValue = -99999.99f; // float

    float ek(time=31, lat=180, lon=360);
      :long_name = "first guess daily product version 1 kriging error per grid";
      :units = "%";
      :code = 23; // int
      :_FillValue = -99999.99f; // float

    float s(time=31, lat=180, lon=360);
      :long_name = "first guess daily product version 1 number of gauges per grid";
      :units = "gauges per gridcell";
      :code = 21; // int
      :_FillValue = -99999.99f; // float

  // global attributes:
  :CDI = "Climate Data Interface version 1.5.9 (http://code.zmaw.de/projects/cdi)";
  :Conventions = "CF-1.4";
  :history = "Fri Feb 05 08:15:42 2016: cdo -setgatts,gattfile gpcc10.nc first_guess_daily_201601.nc\nFri Feb 05 08:15:42 2016: cdo -merge first_guess_daily_precip_201601.nc first_guess_daily_error_201601.nc first_guess_daily_krigingerror_201601.nc first_guess_daily_numgauge_201601.nc gpcc10.nc\nFri Feb 05 08:15:30 2016: cdo cat gpcc10.nc first_guess_daily_numgauge_201601.nc\nFri Feb 05 08:15:30 2016: cdo -b F32 -r -f nc -setgrid,firstguess10desc.asc -settunits,days -setmissval,-99999.99 -invertlatdata -setpartab,codetable.txt -setcode,21 -setdate,2016-01-01 -input,r360x180 gpcc10.nc";
  :DOI = "10.5676/DWD_GPCC/FG_D_100";
  :title = "GPCC first guess daily, version 1.0, precipitation per grid in mm/day, number of gauges per grid, standard deviation per grid in mm/day, kriging error per grid in %, 1.0 degree";
  :summary = "This is the GPCC First Guess Daily Product of daily global land-surface precipitation based on the station database (SYNOP) available via the Global Telecommunication System (GTS) of the World Meteorological Organization (WMO) at the time of analysis (3 - 5 days after end of the analysis month). This product contains the daily totals for a month on a regular latitude/longitude grid with a spatial resolution of 1.0 x 1.0 degree. Interpolation is made for the daily relative quota of the monthly total, i.e., the daily total divided by the monthly total, the latter has the DOI:10.5676/DWD_GPCC/FG_M_100. The temporal coverage of the dataset ranges from January 2009 to the most recent month for which GTS based SYNOP data is available, i.e. the previous month, 3-5 days after its completion.";
  :usage = "This GPCC product is recommended to be used when the timeliness of the precipitation information is of highest importance, e.g. for drought monitoring or climate watch similar to the (monthly) GPCC First Guess Product. In addition the GPCC First Guess Daily product allows to globally study extreme events and related statistics at daily resolution.";
  :keywords = "precipitation climatology,gpcc,global,gpcp,daily";
  :id = "first_guess_daily_precipitation_10";
  :creator_url = "http://gpcc.dwd.de";
  :creator_name = "GPCC/DWD";
  :creator_email = "gpcc@dwd.de";
  :institution = "Deutscher Wetterdienst";
  :date_created = "Fr 5. Feb 08:15:42 UTC 2016";
  :time_coverage_start = "2016-01-01";
  :time_coverage_end = "2016-01-31";
  :time_coverage_resolution = "day";
  :geospatial_lat_min = "-90.";
  :geospatial_lat_max = "90.";
  :geospatial_lon_min = "-180.";
  :geospatial_lon_max = "180.";
  :CDO = "Climate Data Operators version 1.5.9 (http://code.zmaw.de/projects/cdo)";
}